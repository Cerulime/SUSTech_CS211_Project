module Scoreboard(
    input clk, en,
    input [20:0] combo,
    input [1:0] mod,
    input [3:0] difficutly,
    input [20:0] base_score,
    input [20:0] bonus_score,
    input [20:0] acc,
    input [2:0] level,
    output ctr1,
    output [7:0] tube1,
    output ctr2,
    output [7:0] tube2
);

endmodule