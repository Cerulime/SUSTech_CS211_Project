`define NOTE_KEY_BITS 7
`define LENGTH_KEY_BITS 7
`define TUBE_BITS 8
`define CLOCK_BITS 32

`define OCTAVE_BITS 3
`define NOTE_BITS 3
`define LENGTH_BITS 4
`define FULL_NOTE_BITS 3

`define SONG_BITS 3
`define SONG_CNT_BITS 21
`define SCORE_BITS 21
`define REC_CNT_BITS 6