module Controller (
    input clk, rst,
    input [2:0] mode,
    output buzzer
);
endmodule