`define NOTE_KEY_BITS 7
`define LENGTH_KEY_BITS 7
`define TUBE_BITS 8
`define CLOCK_BITS 32

`define OCTAVE_BITS 3
`define NOTE_BITS 3
`define LENGTH_BITS 3
`define FULL_NOTE_BITS 3

`define SONG_BITS 3
`define SONG_CNT_BITS 21
`define SCORE_BITS 21
`define REC_CNT_BITS 6

`define free_mode 1
`define auto_mode 2
`define stdy_mode 3
`define play_mode 4
`define set 5

`define little_star 1
`define two_tigers 2

`define do 0
`define re 1
`define mi 2
`define fa 3
`define so 4
`define la 5
`define xi 6

`define full_note 0
`define half_note 1
`define quarter_note 2
`define eighth_note 3
`define sixteenth_note 4
`define thirty_second_note 5
`define sixty_fourth_note 6

`define zero 8'b11111100
`define one 8'b01100000
`define two 8'b11011010
`define three 8'b11110010
`define four 8'b01100110
`define five 8'b10110110
`define six 8'b10111110
`define seven 8'b11100000
`define eight 8'b11111110
`define nine 8'b11100110
`define A 8'b11101110
`define b 8'b00111110
`define C 8'b10011100
`define c 8'b00011010
`define d 8'b01111010
`define E 8'b10011110
`define F 8'b10001110
`define g 8'b11110110
`define G 8'b10111100
`define H 8'b01101110
`define h 8'b00101110
`define i 8'b10100000
`define I 8'b01100000
`define j 8'b10110000
`define L 8'b00011100
`define l 8'b00001100
`define n 8'b00101010
`define N 8'b11101100
`define O 8'b11111100
`define o 8'b00111010
`define p 8'b11001110
`define q 8'b11100110
`define r 8'b00001010
`define S 8'b10110110
`define t 8'b00011110
`define U 8'b01111100
`define u 8'b00111000
`define y 8'b01110110
`define emp 8'b00000000
