module Seventube(
    input clk, en,
    input float,
    input [22:0] num,
    output ctr1,
    output [7:0] tube1,
    output ctr2,
    output [7:0] tube2
);

endmodule